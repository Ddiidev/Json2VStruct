module type_object

pub enum TypeParser {
	json
	toml
	// yaml
	// xml
	// ini
}
