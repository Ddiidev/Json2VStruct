module entities

pub struct Config {
pub:
	struct_anon                   bool
	omit_empty                    bool = true
	reserved_word_with_underscore bool = true
}
