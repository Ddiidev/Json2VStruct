module contracts

pub interface IGenerator {
	execute(objs KeyValueType) string
}
