module contracts

pub interface INameKey {
mut:
	name string
	attribute_replace_name string
}
