module contracts

pub enum Format {
	json
	yaml
	toml
}
