module contracts

pub struct NameKey {
pub mut:
	name                   string
	attribute_replace_name string
}
