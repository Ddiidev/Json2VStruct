module contracts

pub interface IConfig {
	struct_anon bool
	omit_empty bool
	reserved_word_with_underscore bool
}
