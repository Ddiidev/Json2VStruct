module main

import cli
import os

const str_simple_js = r'
	{
		"name": "André",
		"age": 25
	}
'

fn main() {
	
}
