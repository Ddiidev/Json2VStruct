module entities

pub struct NameKey {
pub mut:
	name       string
	attributes string
}
