module main

const reserved_words = [
	  "if", "is", "else", "for", "in", "fn", "defer", "return", "break",
  "nil", "false", "true", "bool", "int", "float", "string", "rune",
  "i8", "i16", "i32", "i64", "u8", "u16", "u32", "u64", "f32", "f64",
  "char", "voidptr", "any", "type", "struct", "enum", "union", "const",
  "import", "export", "as", "pub", "module", "static", "mut",
  "match"
]
