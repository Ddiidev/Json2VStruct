module parsers

pub enum TypeParser {
	json
	// yaml
	// toml
	// xml
	// ini
}
