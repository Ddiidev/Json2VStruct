module parsers

