module genarators

import contracts

pub struct Generator {
	format contracts.Format
}
