module parsers
