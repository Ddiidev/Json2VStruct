module contracts

pub interface IGenerator {
	execute() string
}
