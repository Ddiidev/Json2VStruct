module main

import x.json2
